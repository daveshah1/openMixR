library ieee ;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--OV16825 Camera Configuration for openMixR 1080p mode

--This configuration is for 1080p, 60fps, 10-bit, 4-lane with a total horizontal length of 4224 pixels
--and a total vertical length of 2496 lines

entity ov16825_1080p_openmixr_regs is
port (clock : in std_logic; --this allows a blockram to be elaborated
  		address : in std_logic_vector(8 downto 0);
  		--This is the I2C data to be written
  		--2 MSBs are address, 1 MSB is data
  		data : out std_logic_vector(23 downto 0));
end ov16825_1080p_openmixr_regs;

architecture behv_cd of ov16825_1080p_openmixr_regs is
begin
	process(clock)
	begin
		if rising_edge(clock) then
			case address(8 downto 0) is
        --Global init
        when "0" & x"00" =>
          data <= x"010301"; --software reset

        when "0" & x"10" => --PLL setup
          data <= x"010000";
        when "0" & x"11" =>
          data <= x"030002";
        when "0" & x"12" =>
          data <= x"030250";
        when "0" & x"13" =>
          data <= x"030501";
        when "0" & x"14" =>
          data <= x"030600";
        when "0" & x"15" =>
          data <= x"030b02";
        when "0" & x"16" =>
          data <= x"030c14";
        when "0" & x"17" =>
          data <= x"030e00";
        when "0" & x"18" =>
          data <= x"031302";
        when "0" & x"19" =>
          data <= x"031414";
        when "0" & x"1a" =>
          data <= x"031f00";

        when "0" & x"20" =>
          data <= x"302201";
        when "0" & x"21" =>
          data <= x"303280";
        when "0" & x"22" =>
          data <= x"3601f8";
        when "0" & x"23" =>
          data <= x"360200";
        when "0" & x"24" =>
          data <= x"360550";
        when "0" & x"25" =>
          data <= x"360600";
        when "0" & x"26" =>
          data <= x"36072b";
        when "0" & x"27" =>
          data <= x"360816";
        when "0" & x"28" =>
          data <= x"360900";
        when "0" & x"29" =>
          data <= x"360e99";
        when "0" & x"2a" =>
          data <= x"360f75";
        when "0" & x"2b" =>
          data <= x"361069";
        when "0" & x"2c" =>
          data <= x"361159";
        when "0" & x"2d" =>
          data <= x"361240";
        when "0" & x"2e" =>
          data <= x"361389";
        when "0" & x"2f" =>
          data <= x"361544";
        when "0" & x"30" =>
          data <= x"361700";
        when "0" & x"31" =>
          data <= x"361820";
        when "0" & x"32" =>
          data <= x"361900";
        when "0" & x"33" =>
          data <= x"361a10";
        when "0" & x"34" =>
          data <= x"361c10";
        when "0" & x"35" =>
          data <= x"361d00";
        when "0" & x"36" =>
          data <= x"361e00";
        when "0" & x"37" =>
          data <= x"364015";
        when "0" & x"38" =>
          data <= x"364154";
        when "0" & x"39" =>
          data <= x"364263";
        when "0" & x"3a" =>
          data <= x"364332";
        when "0" & x"3b" =>
          data <= x"364403";
        when "0" & x"3c" =>
          data <= x"364504";
        when "0" & x"3d" =>
          data <= x"364685";
        when "0" & x"3e" =>
          data <= x"364a07";
        when "0" & x"3f" =>
          data <= x"370708";
        when "0" & x"40" =>
          data <= x"371875";
        when "0" & x"41" =>
          data <= x"371a55";
        when "0" & x"42" =>
          data <= x"371c55";
        when "0" & x"43" =>
          data <= x"373380";
        when "0" & x"44" =>
          data <= x"376000";
        when "0" & x"45" =>
          data <= x"376130";
        when "0" & x"46" =>
          data <= x"376200";
        when "0" & x"47" =>
          data <= x"3763c0";
        when "0" & x"48" =>
          data <= x"376403";
        when "0" & x"49" =>
          data <= x"376500";

        when "0" & x"50" =>
          data <= x"382308";
        when "0" & x"51" =>
          data <= x"382702";
        when "0" & x"52" =>
          data <= x"382800";
        when "0" & x"53" =>
          data <= x"383200";
        when "0" & x"54" =>
          data <= x"383300";
        when "0" & x"55" =>
          data <= x"383400";
        when "0" & x"56" =>
          data <= x"3d8517";
        when "0" & x"57" =>
          data <= x"3d8c70";
        when "0" & x"58" =>
          data <= x"3d8da0";
        when "0" & x"59" =>
          data <= x"3f0002";

        when "0" & x"60" =>
          data <= x"400183";
        when "0" & x"61" =>
          data <= x"400e00";
        when "0" & x"62" =>
          data <= x"401100";
        when "0" & x"63" =>
          data <= x"401200";
        when "0" & x"64" =>
          data <= x"420008";
        when "0" & x"65" =>
          data <= x"43027f";
        when "0" & x"66" =>
          data <= x"4303ff";
        when "0" & x"67" =>
          data <= x"430400";
        when "0" & x"68" =>
          data <= x"430500";
        when "0" & x"69" =>
          data <= x"450130";
        when "0" & x"6a" =>
          data <= x"460320";
        when "0" & x"6b" =>
          data <= x"4b0022";
        when "0" & x"6c" =>
          data <= x"490300";
        when "0" & x"6d" =>
          data <= x"50007f";
        when "0" & x"6e" =>
          data <= x"500101";
        when "0" & x"6f" =>
          data <= x"500400";
        when "0" & x"70" =>
          data <= x"501320";
        when "0" & x"71" =>
          data <= x"505100";
        when "0" & x"72" =>
          data <= x"550001";
        when "0" & x"73" =>
          data <= x"550100";
        when "0" & x"74" =>
          data <= x"550207";
        when "0" & x"75" =>
          data <= x"5503ff";
        when "0" & x"76" =>
          data <= x"55056c";
        when "0" & x"77" =>
          data <= x"550902";
        when "0" & x"78" =>
          data <= x"5780fc";
        when "0" & x"79" =>
          data <= x"5781ff";
        when "0" & x"7a" =>
          data <= x"578740";
        when "0" & x"7b" =>
          data <= x"578808";
        when "0" & x"7c" =>
          data <= x"578a02";
        when "0" & x"7d" =>
          data <= x"578b01";
        when "0" & x"7e" =>
          data <= x"578c01";
        when "0" & x"7f" =>
          data <= x"578e02";
        when "0" & x"80" =>
          data <= x"578f01";
        when "0" & x"81" =>
          data <= x"579001";
        when "0" & x"82" =>
          data <= x"579200";
        when "0" & x"83" =>
          data <= x"598000";
        when "0" & x"84" =>
          data <= x"598121";
        when "0" & x"85" =>
          data <= x"598200";
        when "0" & x"86" =>
          data <= x"598300";
        when "0" & x"87" =>
          data <= x"598400";
        when "0" & x"88" =>
          data <= x"598500";
        when "0" & x"89" =>
          data <= x"598600";
        when "0" & x"8a" =>
          data <= x"598700";
        when "0" & x"8b" =>
          data <= x"598800";

        when "0" & x"90" =>
          data <= x"320115";
        when "0" & x"91" =>
          data <= x"32022a";

        --1080p120 specific config
        when "0" & x"a0" =>
          data <= x"010000";

        when "0" & x"b0" =>
          data <= x"320800";
        when "0" & x"b1" =>
          data <= x"301afb";
        when "0" & x"b2" =>
          data <= x"030264";
        when "0" & x"b3" =>
          data <= x"030501";
        when "0" & x"b4" =>
          data <= x"030e00";
        when "0" & x"b5" =>
          data <= x"30187a";
        when "0" & x"b6" =>
          data <= x"30310a";
        when "0" & x"b7" =>
          data <= x"360305";
        when "0" & x"b8" =>
          data <= x"360402";
        when "0" & x"b9" =>
          data <= x"360a02";
        when "0" & x"ba" =>
          data <= x"360b02";
        when "0" & x"bb" =>
          data <= x"360c12";
        when "0" & x"bc" =>
          data <= x"360d04";
        when "0" & x"bd" =>
          data <= x"361477";
        when "0" & x"be" =>
          data <= x"361631";
        when "0" & x"bf" =>
          data <= x"363140";

        when "0" & x"c0" =>
          data <= x"370060";
        when "0" & x"c1" =>
          data <= x"370110";
        when "0" & x"c2" =>
          data <= x"370222";
        when "0" & x"c3" =>
          data <= x"370340";
        when "0" & x"c4" =>
          data <= x"370410";
        when "0" & x"c5" =>
          data <= x"370501";
        when "0" & x"c6" =>
          data <= x"370604";
        when "0" & x"c7" =>
          data <= x"370840";
        when "0" & x"c8" =>
          data <= x"370978";
        when "0" & x"c9" =>
          data <= x"370a02";
        when "0" & x"ca" =>
          data <= x"370bb2";
        when "0" & x"cb" =>
          data <= x"370c06";
        when "0" & x"cc" =>
          data <= x"370e40";
        when "0" & x"cd" =>
          data <= x"370f0a";

        when "0" & x"d0" =>
          data <= x"371030";
        when "0" & x"d1" =>
          data <= x"371140";
        when "0" & x"d2" =>
          data <= x"371431";
        when "0" & x"d3" =>
          data <= x"371925";
        when "0" & x"d4" =>
          data <= x"371b05";
        when "0" & x"d5" =>
          data <= x"371d05";
        when "0" & x"d6" =>
          data <= x"371e11";
        when "0" & x"d7" =>
          data <= x"371f2d";

        when "0" & x"e0" =>
          data <= x"372015";
        when "0" & x"e1" =>
          data <= x"372130";
        when "0" & x"e2" =>
          data <= x"372215";
        when "0" & x"e3" =>
          data <= x"372330";
        when "0" & x"e4" =>
          data <= x"372408";
        when "0" & x"e5" =>
          data <= x"372508";
        when "0" & x"e6" =>
          data <= x"372604";
        when "0" & x"e7" =>
          data <= x"372704";
        when "0" & x"e8" =>
          data <= x"372804";
        when "0" & x"e9" =>
          data <= x"372904";
        when "0" & x"ea" =>
          data <= x"372a29";
        when "0" & x"eb" =>
          data <= x"372bc9";
        when "0" & x"ec" =>
          data <= x"372ca9";
        when "0" & x"ed" =>
          data <= x"372db9";
        when "0" & x"ee" =>
          data <= x"372e95";
        when "0" & x"ef" =>
          data <= x"372f55";
        when "0" & x"f0" =>
          data <= x"373055";
        when "0" & x"f1" =>
          data <= x"373155";
        when "0" & x"f2" =>
          data <= x"373205";
        when "0" & x"f3" =>
          data <= x"373410";
        when "0" & x"f4" =>
          data <= x"373905";
        when "0" & x"f5" =>
          data <= x"373a40";
        when "0" & x"f6" =>
          data <= x"373b18";
        when "0" & x"f7" =>
          data <= x"373c38";
        when "0" & x"f8" =>
          data <= x"373e15";
        when "0" & x"f9" =>
          data <= x"373f80";

        when "1" & x"00" =>
          data <= x"380001";
        when "1" & x"01" =>
          data <= x"380180";
        when "1" & x"02" =>
          data <= x"380202";
        when "1" & x"03" =>
          data <= x"380394";
        when "1" & x"04" =>
          data <= x"380410";
        when "1" & x"05" =>
          data <= x"3805bf";
        when "1" & x"06" =>
          data <= x"38060b";
        when "1" & x"07" =>
          data <= x"38070f";
        when "1" & x"08" =>
          data <= x"380807";
        when "1" & x"09" =>
          data <= x"380980";
        when "1" & x"0a" =>
          data <= x"380a04";
        when "1" & x"0b" =>
          data <= x"380b38";
        when "1" & x"0c" =>
          data <= x"380c04";
        when "1" & x"0d" =>
          data <= x"380d20";
        when "1" & x"0e" =>
          data <= x"380e09";
        when "1" & x"0f" =>
          data <= x"380fc0";
        when "1" & x"10" =>
          data <= x"381117";
        when "1" & x"11" =>
          data <= x"381302";
        when "1" & x"12" =>
          data <= x"381403";
        when "1" & x"13" =>
          data <= x"381501";
        when "1" & x"14" =>
          data <= x"382000";
        when "1" & x"15" =>
          data <= x"382107";
        when "1" & x"16" =>
          data <= x"382900";
        when "1" & x"17" =>
          data <= x"382a03";
        when "1" & x"18" =>
          data <= x"382b01";
        when "1" & x"19" =>
          data <= x"383008";
        when "1" & x"1a" =>
          data <= x"3f0840";

        when "1" & x"20" =>
          data <= x"400202";
        when "1" & x"21" =>
          data <= x"400304";
        when "1" & x"22" =>
          data <= x"483714";
        when "1" & x"23" =>
          data <= x"350144";
        when "1" & x"24" =>
          data <= x"350808";
        when "1" & x"25" =>
          data <= x"3509ff";
        when "1" & x"26" =>
          data <= x"363800";
        when "1" & x"27" =>
          data <= x"301af0";
        when "1" & x"28" =>
          data <= x"320810";
        when "1" & x"29" =>
          data <= x"3208a0";

        when "1" & x"30" =>
          data <= x"380807";
        when "1" & x"31" =>
          data <= x"380980";
        when "1" & x"32" =>
          data <= x"380a04";
        when "1" & x"33" =>
          data <= x"380b38";
        when "1" & x"34" =>
          data <= x"381000";
        when "1" & x"35" =>
          data <= x"381117";
        when "1" & x"36" =>
          data <= x"381200";
        when "1" & x"37" =>
          data <= x"381302";
        when "1" & x"38" =>
          data <= x"46032f";
        when "1" & x"39" =>
          data <= x"50007f";

        when "1" & x"40" =>
          data <= x"010001";
 				when others =>
						data <= x"000000";
				end case;
		end if;
	end process;
end behv_cd;
